`timescale 1ns / 1ps
//////////////////////////////////////////////////////////////////////////////////
// Company: Boston University
// Engineer: Zafar M. Takhirov
// 
// Create Date:    12:59:40 04/12/2011 
// Design Name: EC311 Support Files
// Module Name:    vga_display 
// Project Name: Lab5 / Lab6 / Project
// Target Devices: xc6slx16-3csg324
// Tool versions: XILINX ISE 13.3
// Description: 
//
// Dependencies: vga_controller_640_60
//
// Revision: 
// Revision 0.01 - File Created
// Additional Comments: 
//
//////////////////////////////////////////////////////////////////////////////////
module vga_display(rst, clk, R, G, B, HS, VS, R_control, G_control, B_control);
    input rst;  // global reset
    input clk;  // 100MHz clk
    
    // color inputs for a given pixel
    input [2:0] R_control, G_control;
    input [1:0] B_control; 
    
    // color outputs to show on display (current pixel)
    output reg [2:0] R, G;
    output reg [1:0] B;
    
    // Synchronization signals
    output HS;
    output VS;
    
    // controls:
    wire [10:0] hcount, vcount; // coordinates for the current pixel
    wire blank; // signal to indicate the current coordinate is blank
    wire figure;    // the figure you want to display
    
    /////////////////////////////////////////////////////
    // Begin clock division
    parameter N = 2;    // parameter for clock division
    reg clk_25Mhz;
    reg [N-1:0] count;
    always @ (posedge clk) begin
        count <= count + 1'b1;
        clk_25Mhz <= count[N-1];
    end
    // End clock division
    /////////////////////////////////////////////////////
    
    // Call driver
    vga_controller_640_60 vc(
        .rst(rst), 
        .pixel_clk(clk_25Mhz), 
        .HS(HS), 
        .VS(VS), 
        .hcounter(hcount), 
        .vcounter(vcount), 
        .blank(blank));
    
    // create a box:
    assign figure = ~blank & (hcount >= 300 & hcount <= 500 & vcount >= 167 & vcount <= 367);

    // send colors:
    always @ (posedge clk) begin
        if (figure) begin   // if you are within the valid region
            R = R_control;
            G = G_control;
            B = B_control;
        end
        else begin  // if you are outside the valid region
            R = 0;
            G = 0;
            B = 0;
        end
    end

endmodule
